<svg x="0" y="0" width="2123.51481" height="1948.03874" version="1.1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink"><g fill="none" stroke="none" stroke-width="2" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10" stroke-dasharray="" stroke-dashoffset="0" font-family="sans-serif" font-weight="normal" font-size="12" text-anchor="start" mix-blend-mode="normal"><line x1="20" y1="203.19393" x2="20" y2="697.26235" stroke="#000000"></line><path d="M20,697.26235c0,0.5 0,0.5 0,0.5c0,7.35035 0.1259,14.761 1.73504,21.93305c1.60914,7.17205 4.68686,14.02759 9.12858,19.88411c4.44173,5.85652 10.16291,10.6664 16.40491,14.54778c6.242,3.88138 12.98463,6.87781 19.71013,9.84352c6.72549,2.96571 13.47235,5.95065 19.72672,9.81208c6.25436,3.86143 11.99693,8.64295 16.47359,14.4728c4.47666,5.82986 7.60307,12.66165 9.26917,19.82069c1.6661,7.15904 1.85623,14.56788 1.92014,21.91795c0.00435,0.49998 0.00435,0.49998 0.00435,0.49998" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="20" y1="697.26235" x2="114.37262" y2="830.49432"></line><polyline points="104.37277,830.54863 114.37262,830.49432 117.74173,821.07895"></polyline></g><line x1="114.37262" y1="830.49432" x2="119.92396" y2="1468.89732" stroke="#000000"></line><path d="M119.92396,1468.89732c0.00435,0.49998 0.00435,0.49998 0.00435,0.49998c0.07191,8.26995 -0.1677,16.53865 -0.60127,24.79754c-0.43357,8.25889 -0.8938,16.65759 1.03169,24.70059c2.33536,9.75507 8.29565,18.4947 16.14292,24.74255c7.84727,6.24785 17.50214,10.0597 27.42786,11.50728c19.85143,2.89517 40.06265,-3.50111 57.64041,-13.1698c17.57777,-9.66869 33.15253,-22.5307 49.62689,-33.97871c16.47436,-11.44801 34.39704,-21.69802 54.17466,-25.06065c16.27595,-2.76727 32.93355,-1.93727 49.41458,-2.90674c0.49914,-0.02936 0.49914,-0.02936 0.49914,-0.02936" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="119.92396" y1="1468.89732" x2="375.28518" y2="1480"></line><polyline points="369.19901,1487.93464 375.28518,1480 369.91065,1471.56707"></polyline></g><line x1="375.28518" y1="1480" x2="752.77565" y2="1457.79464" stroke="#000000"></line><path d="M752.77565,1457.79464c0.49914,-0.02936 0.49914,-0.02936 0.49914,-0.02936c16.47183,-0.96893 32.96508,-1.61293 49.41458,-2.90674c45.4554,-3.57523 91.46422,-14.26524 129.33643,-39.65562c18.93611,-12.69519 35.59319,-28.99827 47.66856,-48.33552c12.07537,-19.33725 19.4654,-41.75504 20.04905,-64.54546c0.42255,-16.49963 -1.78779,-32.94649 -2.6821,-49.42728c-0.02709,-0.49927 -0.02709,-0.49927 -0.02709,-0.49927" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="752.77565" y1="1457.79464" x2="997.03423" y2="1252.39539"></line><polyline points="997.91635,1262.3564 997.03423,1252.39539 987.37223,1249.81745"></polyline></g><line x1="997.03423" y1="1252.39539" x2="958.17491" y2="536.27375" stroke="#000000"></line><path d="M958.17491,536.27375c-0.02709,-0.49927 -0.02709,-0.49927 -0.02709,-0.49927c-0.89412,-16.47728 -2.51164,-32.92664 -2.6821,-49.42728c-0.25879,-25.05073 3.93061,-50.02472 3.06362,-75.06178c-0.43349,-12.51853 -2.15422,-25.07303 -6.23016,-36.91736c-4.07593,-11.84433 -10.58646,-22.98337 -19.72799,-31.54689c-6.02684,-5.64578 -13.03806,-10.11684 -19.99043,-14.57354c-6.95237,-4.4567 -13.83795,-9.01731 -20.61168,-13.74109c-0.41012,-0.28601 -0.41012,-0.28601 -0.41012,-0.28601" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="958.17491" y1="536.27375" x2="891.55896" y2="314.22054"></line><polyline points="901.05317,317.36059 891.55896,314.22054 885.36106,322.06822"></polyline></g><line x1="891.55896" y1="314.22054" x2="469.65777" y2="20" stroke="#000000"></line><path d="M469.65777,20c-0.41012,-0.28601 -0.41012,-0.28601 -0.41012,-0.28601c-6.79695,-4.73997 -13.34872,-9.81903 -19.73515,-15.09912c-6.38643,-5.28009 -12.96376,-10.72449 -20.86696,-13.21551c-4.9239,-1.55197 -10.22129,-1.83823 -15.31362,-0.98877c-5.09233,0.84947 -9.9775,2.8213 -14.32499,5.60568c-8.69497,5.56877 -15.09554,14.2833 -19.03351,23.82826c-7.87593,19.08991 -6.23347,40.55002 -5.55017,61.1895c0.54597,16.49116 0.56887,32.9949 0.85331,49.49264c0.00862,0.49993 0.00862,0.49993 0.00862,0.49993" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="469.65777" y1="20" x2="375.28518" y2="131.02661"></line><polyline points="372.75849,121.35108 375.28518,131.02661 385.24138,131.96153"></polyline></g><line x1="375.28518" y1="131.02661" x2="380.83646" y2="453.00378" stroke="#000000"></line><path d="M380.83646,453.00378c0.00862,0.49993 0.00862,0.49993 0.00862,0.49993c0.14262,8.27204 -0.04865,16.54529 -0.44776,24.80892c-0.39911,8.26364 -0.82357,16.68792 1.30107,24.68372c2.5934,9.75992 9.13481,18.32667 17.62549,23.79385c8.49068,5.46718 18.82498,7.87393 28.90043,7.19043c10.07544,-0.6835 19.864,-4.38807 28.15078,-10.15963c8.28678,-5.77156 15.08963,-13.5651 20.11621,-22.32382c10.05316,-17.51744 12.87601,-38.43542 11.5782,-58.59087c-1.29781,-20.15546 -6.47096,-39.83258 -11.52359,-59.38757c-5.05264,-19.55499 -10.0347,-39.30149 -10.93613,-59.47856c-0.90143,-20.17707 2.5527,-41.05841 13.28654,-58.16722c5.36692,-8.55441 12.51545,-16.04727 21.07572,-21.40483c8.56027,-5.35756 18.54746,-8.53155 28.64567,-8.6201c10.09821,-0.08855 20.27261,2.97792 28.3674,9.01581c8.09478,6.03789 13.99692,15.07833 15.81576,25.01179c1.49018,8.13855 0.37287,16.50386 -0.70581,24.7071c-1.07867,8.20324 -1.94843,16.43351 -2.48112,24.6902c-0.03219,0.49896 -0.03219,0.49896 -0.03219,0.49896" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="380.83646" y1="453.00378" x2="569.58176" y2="319.77187"></line><polyline points="569.61973,329.7718 569.58176,319.77187 560.17191,316.38738"></polyline></g><line x1="569.58176" y1="319.77187" x2="547.3764" y2="663.95437" stroke="#000000"></line><path d="M547.3764,663.95437c-0.03219,0.49896 -0.03219,0.49896 -0.03219,0.49896c-0.53272,8.25713 -1.40563,16.48756 -2.48936,24.69058c-1.08374,8.20302 -2.20631,16.57114 -0.69756,24.70672c1.84315,9.93876 7.81269,18.9598 15.96277,24.93911c8.15009,5.97931 18.36399,8.95285 28.47067,8.77674c10.10668,-0.17611 20.07321,-3.42888 28.6175,-8.82991c8.54429,-5.40103 15.68403,-12.90216 21.09533,-21.43995c10.82261,-17.07558 14.59498,-37.83106 14.44995,-58.04697c-0.14503,-20.21592 -3.95822,-40.19814 -7.23633,-60.14704c-3.27813,-19.94889 -6.03885,-40.21391 -4.06445,-60.33371c1.97439,-20.1198 9.0985,-40.31748 23.24272,-54.76204c7.07211,-7.22228 15.82166,-12.87578 25.47476,-15.87475c9.6531,-2.99897 20.20776,-3.27901 29.87178,-0.31542c9.66402,2.96359 18.36328,9.23689 23.82111,17.74503c5.45782,8.50813 7.52592,19.22767 5.1565,29.05426c-1.94032,8.04697 -6.53641,15.16025 -11.01693,22.12039c-4.48052,6.96014 -8.7703,14.04246 -12.74364,21.30408c-0.24001,0.43863 -0.24001,0.43863 -0.24001,0.43863" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="547.3764" y1="663.95437" x2="725.01902" y2="558.47911"></line><polyline points="724.26918,568.45095 725.01902,558.47911 715.90501,554.36392"></polyline></g><line x1="564.03042" y1="852.69955" x2="725.01902" y2="558.47911" stroke="#000000"></line><path d="M564.03042,852.69955c-0.24001,0.43863 -0.24001,0.43863 -0.24001,0.43863c-3.96839,7.25256 -8.18739,14.36415 -12.55877,21.38119c-4.37138,7.01704 -8.82378,14.12541 -11.2018,22.04329c-2.87467,9.57151 -2.43675,19.95251 0.20722,29.5903c2.64397,9.63779 7.41487,18.58638 13.06035,26.83296c11.29096,16.49316 26.09487,30.37531 37.12471,47.04423c5.51492,8.33446 10.0783,17.4055 12.41746,27.12176c2.33917,9.71627 2.36679,20.12833 -0.95669,29.5534c-3.32348,9.42507 -10.17888,17.75855 -19.26474,21.92083c-4.54293,2.08114 -9.5841,3.1039 -14.57302,2.82101c-4.98892,-0.28288 -9.91458,-1.88537 -14.03987,-4.70519c-6.85244,-4.68394 -11.15084,-12.18478 -15.26536,-19.39351c-4.11452,-7.20873 -8.4938,-14.26531 -13.28045,-21.0464c-0.28834,-0.40848 -0.28834,-0.40848 -0.28834,-0.40848" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="564.03042" y1="852.69955" x2="525.1711" y2="1035.89357"></line><polyline points="518.34807,1028.58288 525.1711,1035.89357 534.37452,1031.98242"></polyline></g><line x1="525.1711" y1="1035.89357" x2="325.32318" y2="752.77568" stroke="#000000"></line></g></svg>