<svg x="0" y="0" width="1868.10278" height="1326.50995" version="1.1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink"><g fill="none" stroke="none" stroke-width="2" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10" stroke-dasharray="" stroke-dashoffset="0" font-family="sans-serif" font-weight="normal" font-size="12" text-anchor="start" mix-blend-mode="normal"><polyline points="284.8006,662.23563 274.46392,662.56109 263.58345,662.7457 252.32883,662.79942 240.86965,662.73208 229.37555,662.55352 218.01614,662.27357 206.9611,661.90207 196.38003,661.44886 186.44252,660.92376 177.31828,660.33662" stroke="#000000"></polyline><polyline points="185.08607,666.0891 185.28684,661.71432 185.57717,657.01517 186.02914,652.09162 186.71475,647.04356 187.70614,641.97107 189.07529,636.97402 190.89437,632.15218 193.23541,627.60576 196.17045,623.43451 199.77159,619.73842 204.37524,616.08826 208.72587,613.24564 212.90036,611.02539 216.97568,609.2429 221.02862,607.71345 225.13621,606.25198 229.37523,604.67378 233.82264,602.79406 238.55536,600.42806 243.65023,597.39082 245.51232,595.6908 247.30162,593.03782 248.99516,589.42777 250.57017,584.85637 252.00364,579.31959 253.27271,572.81319 254.35446,565.33308 255.22609,556.87503 255.86457,547.435 256.24704,537.00877 256.60206,527.87377 257.14801,519.18068 257.74283,510.83845 258.24441,502.75586 258.51063,494.84177 258.39946,487.00496 257.76877,479.15427 256.4764,471.19851 254.3804,463.04657 251.33852,454.60723 247.31908,445.21778 243.47804,436.70715 239.86048,428.86635 236.51157,421.48638 233.47638,414.3582 230.80005,407.27288 228.52765,400.02138 226.7043,392.39464 225.37519,384.18374 224.58528,375.17963 224.3998,370.93812 224.33138,365.87747 224.4993,360.00144 225.02266,353.31389 226.02064,345.81859 227.61241,337.51944 229.91719,328.42016 233.05408,318.52459 237.14232,307.83656 242.30096,296.35987" stroke="#000000"></polyline><path d="M185.08607,666.0891c-0.01375,0.29968 -0.01375,0.29968 -0.01375,0.29968c-0.22724,4.95154 -0.31536,9.90815 -0.31659,14.8649c-0.00123,4.95675 0.01004,9.96071 -1.04502,14.80387c-1.25061,5.74082 -4.06501,11.13439 -8.06654,15.43658c-4.00152,4.30219 -9.18017,7.50044 -14.82178,9.14158c-5.6416,1.64114 -11.7307,1.71938 -17.40988,0.2134c-5.67918,-1.50597 -10.93175,-4.59305 -15.00284,-8.82947c-4.07109,-4.23642 -6.9477,-9.61055 -8.20475,-15.34996c-1.25706,-5.73941 -0.88945,-11.82692 1.05918,-17.36984c1.94863,-5.54291 5.47343,-10.52345 10.05944,-14.19626c4.58601,-3.67281 10.21934,-6.02503 16.05666,-6.69345c4.92536,-0.564 9.90255,0.01089 14.82877,0.56731c4.92622,0.55642 9.86261,1.02156 14.80993,1.33992c0.29938,0.01926 0.29938,0.01926 0.29938,0.01926" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="185.08607" y1="666.0891" x2="177.31828" y2="660.33662"></line><polyline points="186.80273,657.16722 177.31828,660.33662 177.05267,670.3331"></polyline></g><polyline points="217.03269,160.40316 216.84473,181.21314 215.09883,198.97465 212.02587,214.20909 207.85683,227.43801 202.82266,239.18292 197.15422,249.96536 191.08255,260.3068 184.8386,270.7287 178.65317,281.75267 172.75737,293.9001 171.81364,298.57207 170.76832,304.74863 169.77353,312.23653 168.9814,320.84249 168.54413,330.37326 168.61379,340.63547 169.34268,351.43601 170.88289,362.58147 173.3866,373.87862 177.00601,385.13422 179.25576,390.28626 182.49702,396.26248 186.78554,402.89297 192.17717,410.00774 198.72761,417.43705 206.49265,425.01093 215.52815,432.55946 225.88986,439.91279 237.63353,446.90099 250.81499,453.35426" stroke="#000000"></polyline><path d="M250.81499,453.35426c0.26944,0.13191 0.26944,0.13191 0.26944,0.13191c3.22273,1.57775 6.48126,3.12219 9.92423,4.13274c3.44297,1.01055 7.04847,1.48398 10.63288,1.31897c7.16883,-0.33001 13.92579,-3.2801 20.37783,-6.42212c6.45204,-3.14202 13.08494,-6.28814 20.22586,-7.00118c3.57046,-0.35652 7.19395,-0.11707 10.70006,0.64612c3.50611,0.76319 6.87329,2.04966 10.20897,3.372c0.27889,0.11056 0.27889,0.11056 0.27889,0.11056" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="250.81499" y1="453.35426" x2="333.43315" y2="449.64325"></line><polyline points="328.07073,458.0839 333.43315,449.64325 327.33559,441.71736"></polyline></g><polyline points="333.43315,449.64325 346.84981,454.96192 358.84619,460.47574 370.02234,466.01647 380.9781,471.41577 392.31336,476.5055 404.62817,481.11732 418.52232,485.08298 434.59585,488.23425 453.44857,490.40289 475.68051,491.42054 487.81314,491.07077 502.05425,489.53126 518.51323,486.60017 537.29953,482.07596 558.52263,475.75688 582.29192,467.44119 608.71684,456.92724 637.90688,444.01329 669.97138,428.49776 705.01977,410.17884" stroke="#000000"></polyline><path d="M705.01977,410.17884c0.26587,-0.13897 0.26587,-0.13897 0.26587,-0.13897c4.41077,-2.3054 8.9459,-4.3615 13.54743,-6.25774c4.60153,-1.89623 9.37273,-3.86652 12.77403,-7.49983c3.15264,-3.3677 4.80163,-8.04162 4.68658,-12.65327c-0.11505,-4.61165 -1.94448,-9.12451 -4.89905,-12.66726c-2.95457,-3.54275 -6.99515,-6.1247 -11.38453,-7.5438c-4.38938,-1.41911 -9.11429,-1.69734 -13.68023,-1.03951c-9.13188,1.31565 -17.41181,6.27658 -24.26798,12.45033c-6.85617,6.17374 -12.48091,13.56444 -18.25727,20.75859c-5.77636,7.19416 -11.82484,14.31074 -19.29775,19.72164c-7.47291,5.4109 -16.58493,9.03236 -25.78872,8.39015c-4.6019,-0.3211 -9.15377,-1.72097 -13.01589,-4.24379c-3.86212,-2.52282 -7.0087,-6.18788 -8.7026,-10.47872c-1.6939,-4.29084 -1.88615,-9.19816 -0.31572,-13.53571c1.57043,-4.33755 4.93835,-8.03815 9.2,-9.8042c4.60111,-1.90672 9.78145,-1.59286 14.75232,-1.28252c4.97087,0.31034 9.95266,0.4367 14.93029,0.26629c0.29982,-0.01026 0.29982,-0.01026 0.29982,-0.01026" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="705.01977" y1="410.17884" x2="635.86638" y2="384.61026"></line><polyline points="644.08695,378.9162 635.86638,384.61026 638.40544,394.28255"></polyline></g><polyline points="635.86638,384.61026 648.80102,384.16742 660.37959,384.86562 670.80939,386.79235 680.29795,390.03517 689.05259,394.68153 697.28073,400.81896 705.19001,408.53503 712.98752,417.91718 720.88102,429.05291 729.0776,442.02981 733.71061,449.05687 739.27209,456.44852 745.63365,464.14816 752.66633,472.09943 760.2415,480.24575 768.23045,488.53069 776.50452,496.89761 784.9349,505.29016 793.39283,513.65179 801.74971,521.92603 809.42714,530.37115 815.78837,539.01111 820.87881,547.69674 824.74341,556.27903 827.42757,564.60894 828.97627,572.53746 829.43467,579.91548 828.84807,586.59395 827.26155,592.42388 824.72028,597.25614 822.44047,599.90204 819.80408,601.95757 816.83164,603.56187 813.54348,604.85407 809.96001,605.97355 806.10179,607.05919 801.98923,608.25043 797.64277,609.68639 793.08284,611.50617 788.32985,613.84899 785.0124,616.16112 781.80216,619.35125 778.77103,623.29648 775.99089,627.87404 773.5336,632.96101 771.47094,638.4344 769.8748,644.17153 768.81693,650.04939 768.36934,655.9452 768.60368,661.73594" stroke="#000000"></polyline><path d="M768.60368,661.73594c0.01213,0.29975 0.01213,0.29975 0.01213,0.29975c0.20056,4.95597 0.5706,9.90312 1.04602,14.84031c0.47542,4.93719 0.96986,9.94278 0.15488,14.8354c-0.80876,4.85529 -2.96729,9.47857 -6.17021,13.21611c-3.20293,3.73754 -7.44106,6.57863 -12.11513,8.1217c-4.67406,1.54307 -9.77066,1.78371 -14.56935,0.68804c-4.79869,-1.09567 -9.28574,-3.52449 -12.82707,-6.9431c-3.54133,-3.41861 -6.12683,-7.8172 -7.39127,-12.57421c-1.26444,-4.75701 -1.20424,-9.85881 0.17198,-14.58469c1.37622,-4.72588 4.06449,-9.06233 7.68503,-12.39694c3.62054,-3.33461 8.16297,-5.65787 12.98581,-6.64182c4.8599,-0.99151 9.88004,-0.6797 14.83125,-0.3844c4.95121,0.2953 9.90854,0.48502 14.86851,0.5052c0.3,0.00122 0.3,0.00122 0.3,0.00122" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="768.60368" y1="661.73594" x2="767.58624" y2="660.7185"></line><polyline points="777.43431,658.98202 767.58624,660.7185 765.84976,670.56658"></polyline></g><polyline points="767.58624,660.7185 776.43578,660.75449 784.99889,660.79362 793.48774,660.83091 802.11429,660.86139 811.09073,660.8802 820.6289,660.88236 830.94099,660.86291 842.23896,660.81686 854.73498,660.73936 868.64091,660.62533" stroke="#000000"></polyline><path d="M868.64091,660.62533c0.29999,-0.00246 0.29999,-0.00246 0.29999,-0.00246c9.89971,-0.08118 19.80056,-0.06557 29.699,-0.24354c26.73416,-0.48069 53.68993,-2.89709 79.16564,-11.01709c25.47571,-8.12 49.53978,-22.29971 66.19032,-43.22113c8.32527,-10.46071 14.70931,-22.52183 18.20958,-35.42472c3.50027,-12.90289 4.07651,-26.64728 1.19457,-39.7022c-2.88194,-13.05492 -9.26765,-25.38371 -18.61569,-34.94147c-9.34804,-9.55776 -21.67266,-16.26193 -34.86122,-18.45247c-9.77026,-1.62278 -19.74516,-1.41633 -29.62389,-2.12494c-0.29923,-0.02146 -0.29923,-0.02146 -0.29923,-0.02146" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="868.64091" y1="660.62533" x2="980" y2="475.47385"></line><polyline points="984.06342,484.61106 980,475.47385 970.02406,476.1671"></polyline></g><polyline points="980,475.47385 964.69476,474.37599 951.49767,470.41822 940.25991,464.05034 930.83242,455.72216 923.06625,445.88339 916.81256,434.98389 911.92231,423.47348 908.24654,411.8019 905.63641,400.41898 903.94288,389.77446 902.52465,376.89548 901.37599,363.4966 900.37563,349.76885 899.40251,335.90335 898.33557,322.09103 897.05363,308.52298 895.43555,295.39026 893.36024,282.88381 890.70667,271.19478 887.35354,260.51411 886.14771,258.18637 884.57631,255.22014 882.49312,251.89658 879.75167,248.4966 876.2056,245.30123 871.70868,242.59155 866.11445,240.6485 859.27654,239.75314 851.04862,240.18653 841.28432,242.22962" stroke="#000000"></polyline><path d="M841.28432,242.22962c-0.29364,0.06144 -0.29364,0.06144 -0.29364,0.06144c-4.85047,1.01492 -9.72564,1.90651 -14.61382,2.72066c-4.88818,0.81415 -9.8164,1.62269 -14.45662,3.36207c-7.48863,2.8071 -13.96615,8.10093 -18.50166,14.68793c-4.53552,6.587 -7.1545,14.42416 -7.84621,22.39165c-1.38342,15.93499 4.91466,31.88635 14.82168,44.44376c9.90702,12.55741 23.19146,22.04987 37.07789,29.98741c13.88644,7.93754 28.52667,14.48213 42.5117,22.24465c13.98503,7.76251 27.47551,16.89439 37.84851,29.06971c10.373,12.17532 17.44129,27.72184 17.06057,43.71223c-0.19036,7.9952 -2.2587,15.98231 -6.28546,22.89205c-4.02676,6.90975 -10.0401,12.70415 -17.25335,16.1579c-7.21325,3.45375 -15.61583,4.49695 -23.37872,2.57422c-7.76289,-1.92273 -14.79834,-6.86727 -18.95055,-13.70237c-2.57458,-4.2381 -4.05121,-9.03642 -5.52162,-13.77222c-1.47041,-4.7358 -3.0356,-9.442 -4.7507,-14.09478c-0.10376,-0.28148 -0.10376,-0.28148 -0.10376,-0.28148" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="841.28432" y1="242.22962" x2="858.64855" y2="454.68445"></line><polyline points="850.01702,449.63503 858.64855,454.68445 866.34561,448.30047"></polyline></g><polyline points="858.64855,454.68445 853.82671,441.60367 849.82505,429.00632 846.60758,416.75177 844.13873,404.69945 842.38239,392.70869 841.30302,380.63892 840.86472,368.34951 841.03172,355.69995 841.76823,342.54951 843.03849,328.75772 844.50147,313.06806 845.40185,297.82426 845.63673,283.13836 845.10277,269.12234 843.69708,255.8884 841.31642,243.54841 837.8578,232.2145 833.21821,221.99877 827.29441,213.01315 819.9834,205.36977 797.43005,189.63622 773.86154,180.25791 748.28106,176.0551 719.69237,175.84816 687.099,178.45737 649.50436,182.70309 605.91204,187.40554 555.32558,191.38504 496.74856,193.46196 429.18445,192.45658" stroke="#000000"></polyline><path d="M429.18445,192.45658c-0.29997,-0.00446 -0.29997,-0.00446 -0.29997,-0.00446c-9.89915,-0.1473 -19.79678,-0.52173 -29.69671,-0.4419c-28.71828,0.23156 -57.66735,5.708 -83.41795,18.42413c-25.7506,12.71613 -48.16011,32.95899 -61.16957,58.56265c-4.48507,8.82698 -8.11709,18.05852 -12.1763,27.08925c-0.12299,0.27363 -0.12299,0.27363 -0.12299,0.27363" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="429.18445" y1="192.45658" x2="242.30096" y2="296.35987"></line><polyline points="243.33354,286.41333 242.30096,296.35987 251.29449,300.73211"></polyline></g><polyline points="340.81511,255.17669 335.50407,267.82236 332.80277,279.7674 332.49721,290.93723 334.37336,301.25748 338.2172,310.65346 343.81468,319.05087 350.95188,326.37501 359.41479,332.55152 368.98929,337.50576 379.46146,341.16332" stroke="#000000"></polyline><path d="M379.46146,341.16332c0.28322,0.09892 0.28322,0.09892 0.28322,0.09892c4.67894,1.63419 9.40041,3.14297 14.14583,4.57265c4.74542,1.42968 9.53532,2.85986 13.89318,5.22039c5.92758,3.21081 10.88505,8.1866 14.07213,14.12698c3.18708,5.94037 4.5915,12.82307 3.9845,19.53701c-0.607,6.71395 -3.2234,13.23369 -7.42764,18.5034c-4.20424,5.26971 -9.98057,9.26916 -16.39333,11.3481c-6.41276,2.07894 -13.43756,2.22914 -19.93277,0.42421c-6.49521,-1.80493 -12.43583,-5.55835 -16.85329,-10.65066c-4.41746,-5.09231 -7.2945,-11.50406 -8.15976,-18.18963c-0.86526,-6.68557 0.28491,-13.61911 3.26435,-19.66629c2.19049,-4.44588 5.27915,-8.37749 8.33127,-12.28244c3.05212,-3.90495 6.03847,-7.86117 8.91675,-11.89597c0.17422,-0.24423 0.17422,-0.24423 0.17422,-0.24423" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="379.46146" y1="341.16332" x2="377.76014" y2="342.06575"></line><polyline points="378.98872,332.14151 377.76014,342.06575 386.66568,346.61453"></polyline></g><polyline points="377.76014,342.06575 381.24,337.18766 383.61725,332.58622 385.17826,328.10194 386.20954,323.57552 386.9974,318.84745 387.82827,313.75831 388.9886,308.14872 390.76477,301.85921 393.44326,294.73033 397.3104,286.60277 400.79583,280.62368 404.96562,274.26623 409.54134,267.46913 414.24449,260.17104 418.7967,252.31067 422.91947,243.82674 426.33431,234.65795 428.7628,224.74298 429.92642,214.02059 429.54676,202.42943 427.69115,188.02819 425.0854,174.85753 421.4773,162.51894 416.61466,150.614 410.24532,138.74425 402.11711,126.51123 391.9778,113.51649 379.57522,99.36155 364.65715,83.64798 346.97141,65.97729 331.12362,52.18299 315.05483,41.37953 298.84759,33.22108 282.58441,27.36181 266.34798,23.45592 250.22072,21.15752 234.28532,20.12084 218.6243,20 203.32024,20.44919 188.45568,21.12258 178.47558,22.36995 168.35897,25.15259 158.01221,29.39879 147.3417,35.037 136.25378,41.99553 124.65481,50.20275 112.45114,59.58709 99.54917,70.07685 85.85523,81.60042 71.27569,94.08618 68.52281,96.78788 66.62796,99.34931 65.42566,101.8046 64.75032,104.18793 64.43649,106.5334 64.31856,108.87522 64.23106,111.24752 64.00848,113.68443 63.48525,116.22011 62.49586,118.88874 58.83485,125.69886 54.23443,132.78918 48.99781,140.07803 43.42827,147.48375 37.82898,154.92474 32.50324,162.31935 27.75423,169.58588 23.88519,176.64272 21.19938,183.40821 20,189.80073 20.32367,194.19572 21.68135,198.6239 23.89868,203.07586 26.80134,207.54208 30.215,212.013 33.9653,216.47923 37.87789,220.93118 41.77846,225.35941 45.49268,229.7544 48.84619,234.10665 51.13307,237.52641 53.46292,241.37745 55.85187,245.51189 58.3161,249.78193 60.8717,254.03971 63.53484,258.13735 66.32163,261.92694 69.24824,265.26066 72.3308,267.99066 75.58543,269.969 80.95449,271.52732 87.34901,271.84748 94.56793,271.06691 102.41011,269.32312 110.67446,266.75358 119.15991,263.49574 127.66535,259.68718 135.98963,255.46524 143.93172,250.9675 151.2905,246.33142" stroke="#000000"></polyline><path d="M151.2905,246.33142c0.25383,-0.15991 0.25383,-0.15991 0.25383,-0.15991c4.21605,-2.65614 8.59107,-5.04783 13.05194,-7.26838c2.23044,-1.11027 4.46182,-2.23259 6.55141,-3.5895c2.08958,-1.3569 4.04583,-2.96894 5.5255,-4.97347c2.29842,-3.11372 3.3259,-7.08212 3.11444,-10.94648c-0.21146,-3.86436 -1.61697,-7.61683 -3.75566,-10.84235c-4.27739,-6.45104 -11.23033,-10.64339 -18.35121,-13.67735c-7.12089,-3.03396 -14.63643,-5.12974 -21.57522,-8.55977c-3.4694,-1.71501 -6.79273,-3.76847 -9.68483,-6.34019c-2.8921,-2.57172 -5.34829,-5.67773 -6.91408,-9.21698c-2.00841,-4.53974 -2.53533,-9.57481 -3.06217,-14.51094c-0.52683,-4.93613 -1.17866,-9.85865 -2.02974,-14.74932c-0.05143,-0.29556 -0.05143,-0.29556 -0.05143,-0.29556" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="151.2905" y1="246.33142" x2="114.36326" y2="141.20124"></line><polyline points="123.99272,143.89817 114.36326,141.20124 108.53549,149.32756"></polyline></g><polyline points="207.41734,73.86495 210.28996,72.04231 213.52992,70.70752 217.04696,69.838 220.75078,69.41116 224.55107,69.40443 228.35763,69.79525 232.08015,70.56106 235.62832,71.67926 238.91189,73.12733 241.84055,74.88266 244.52785,76.9972 246.93147,79.58049 249.03828,82.59441 250.83526,86.00088 252.30926,89.76182 253.44717,93.83911 254.23594,98.19465 254.66241,102.79039 254.71353,107.58821 254.37613,112.54999" stroke="#000000"></polyline><path d="M254.37613,112.54999c-0.02035,0.29931 -0.02035,0.29931 -0.02035,0.29931c-0.34734,5.10804 0.0149,10.23044 0.7996,15.28979c0.39235,2.52967 0.75923,5.09609 0.49084,7.6419c-0.13419,1.27291 -0.43398,2.5355 -0.97169,3.69704c-0.53771,1.16154 -1.32023,2.22104 -2.33369,3.00284c-1.35364,1.04422 -3.08008,1.55417 -4.78965,1.56372c-1.70957,0.00954 -3.40146,-0.46187 -4.93474,-1.21803c-3.06657,-1.51231 -5.45268,-4.08697 -7.77927,-6.59255c-2.32659,-2.50557 -4.74738,-5.0573 -7.84711,-6.50041c-1.54987,-0.72156 -3.25649,-1.14575 -4.96477,-1.07868c-1.70828,0.06707 -3.41623,0.64556 -4.72165,1.74946c-0.97844,0.82739 -1.70924,1.92641 -2.18559,3.11595c-0.47635,1.18954 -0.7055,2.46889 -0.76575,3.74885c-0.1205,2.55991 0.40544,5.10253 0.95509,7.60564c1.09929,5.00622 1.77429,10.10306 1.728,15.22834c-0.00271,0.29999 -0.00271,0.29999 -0.00271,0.29999" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="254.37613" y1="112.54999" x2="217.03269" y2="160.40316"></line><polyline points="214.10357,150.84177 217.03269,160.40316 227.01928,160.92087"></polyline></g><polyline points="114.36326,141.20124 114.33299,141.02732 114.27008,140.53555 114.21626,139.77085 114.21328,138.77813 114.30292,137.60237 114.52693,136.28847 114.92707,134.88137 115.54513,133.42601 116.4228,131.96736 117.60192,130.55029 119.01528,129.28603 120.52882,128.24211 122.08392,127.39799 123.62191,126.73311 125.08416,126.22693 126.41203,125.85886 127.54691,125.60837 128.43013,125.45488 129.00305,125.37787 129.20707,125.35676" stroke="#000000"></polyline><path d="M129.20707,125.35676c0.29841,-0.03087 0.29841,-0.03087 0.29841,-0.03087c7.91983,-0.81926 15.91372,-2.06998 23.12835,-5.43807c7.21462,-3.36809 13.43392,-8.55959 18.98659,-14.26596c5.55267,-5.70637 10.65729,-11.85034 16.45796,-17.30443c5.80066,-5.45409 12.36265,-10.02608 19.08566,-14.29176c0.25331,-0.16072 0.25331,-0.16072 0.25331,-0.16072" stroke="#ff0000"></path><g stroke="#ff0000"><line x1="129.20707" y1="125.35676" x2="207.41734" y2="73.86495"></line><polyline points="207.13114,83.86086 207.41734,73.86495 198.12215,70.17721"></polyline></g></g></svg>